
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:  Fudan University
// Engineer: Gu Chenghao, Ye HanChen, Zhang Bingyi
// 
// Create Date: 11/17/2017 08:42:11 AM
// Design Name: 
// Module Name: simulate_163length_4digital
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module simulate_163length_4digital;


parameter DATA_WIDTH = 163;
parameter DIGITAL = 4;
parameter ITN = 41;
parameter DATA_WIDTH_BIN = 164;

reg rst;
reg clk;
reg start;
reg [DATA_WIDTH - 1 : 0] a;
reg [DATA_WIDTH - 1 : 0] g;
reg [DIGITAL - 1:0] b;
	
wire [DATA_WIDTH - 1 : 0] t_i_j;
wire done;

gf2m inst_gf2m
(
	.rst(rst),
	.clk(clk),
	.start(start),
	.a(a),
	.g(g),
	.b(b),
	
	.t_i_j(t_i_j),
	.done(done)
);


reg [DATA_WIDTH_BIN - 1 : 0] b_total;
reg [DATA_WIDTH - 1 : 0] t_expected;

always
begin
    clk = 1'b0;
    #10;
    clk = 1'b1;
    #10;
end

initial begin
// initial state
a = 163'd0;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'd0;
t_expected = 163'd0;
rst = 1'b0;
start = 1'b0;
#100;
rst = 1'b1;
#100;

start = 1'b1;
a = 163'b1101100110001101100111001110110001001101000010100000000011111001110111100000110001001100011100001011001010000001110101000011000001111001000011101100011110010000010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00111111111111111010011111010100011111110000101111111100111100110011101001110010111110000000100110101110011101111000001010101101011000100011111000110100110100111000;
t_expected = 163'b1101100000000011010001111000000011001110110001100011010000110011011010011101111100000011001000111100011111110010010010111111000000000111101010010011000101010100100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0111001100101100111000110010001111111011010111101001100000111101011010100110000111110010110101101101101010101010010011001111010110010101111011111000110010001010100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01010100101011101110000010011011011011001011011101010001110110100001000100111011001001101100000101000110100111001110101100100100110100000110001101101110000001111011;
t_expected = 163'b0101110001110001110101000111011000100111010000110111000101001000011010001111001110001011001000101100111111111011101000110001010000110101010000011011110011111010111;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0100010111010101000101110111111011011010010110011100010101100111000001110000110001111000000110110001101110100010111100100011101001010100100100111110100100110000110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00001110010100000000101010111011010011011000001100110011000010010001010111110010110101010110100000011101101001010111100011011001011101000111110010100001011110111111;
t_expected = 163'b0101100110001101001010000100011001000111100101001001011011110110001100001001101111010010011010110011011001101111011000010111001000000111100100000011110000011100010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0101111101100101110000001001000011100110110110010100011110100100011010100100100111000011111111101101010011001101100100001010000100101000010110111000011010110011000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01110101001100001000110100100111111111000001101110101010011110001011111000010011000100100111000000000001000011100011001111010001010000100011101111111110001001101100;
t_expected = 163'b0000001001101111111101101110110001101010111111000000001100011111001111101011000110100001100110011001011110010100000111111110000010000100011110011000001010011101001;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1111001101001000101000110101011101000000100011010101111000001110000101110011000101011001010110011010010011110101001010000110111011000010101100111110100000101001110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01001111011000010100111100000101111111110110011110000011011110001101110100011011111011001101101101001010001001010111000000001000101100011110010000011000110010101101;
t_expected = 163'b1110110010000111101001011111101001000100110101010111000001110010111000101101001010011110000011011110011101000111011001010011111110101011000111001010111100011001010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1100000111111001010101010000101001111100000010011100011001000110011110100101110011110011100011000110111111110111100110101010111000000110010110100001101100000011100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00010100000110011011000000010101110001101101011101010001000010011101000111011010001011111101001010110011111111001010100110010001001101111011000100000011100101111111;
t_expected = 163'b0100100110001100110000110110100110001110111001100001011001110100000011111101110010100100110001100100001001001001000000011011100000111111100000001010111000000101100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1110111101000000111000001100010001011111000001100111111010010000000000110001100101101001001010000010101010011110011001000100000111111111010100100111010010010001010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01111110011110010011011111111011111001101110101101111000110010000111101010100111110110000010001011101011010101111100101011011101000000011111111011001100011010110000;
t_expected = 163'b0111110101100010101100111110111001010000011101000010110011000010101111100011000101101010100000011001110101010011110000011100001011001001010001000110010111110110110;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0101011110010000101111110000000111100011110000100010001111011011101001100111010001010000110011111110001010010110110001011101101000011011101111100001001100001011000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01000101101001001101110111111011111001111101010110011000111100110011101101101110010001111010101111100100011011000000000101100100101100111110100110001010000101110001;
t_expected = 163'b1101110101101010100010111111000011100100001101001010100000111100111110110111101001110101000001101000011110010110100101010000110101100010110001010110011000110111100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0100000010111001010110010110111111000111110100101011101100011011110010110001000111001010111010100000000111111100011111111001011110010001010011100101100001100000100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00111111110101000001101011001111110101000110010110000011101000100001010111101110101000011000001110011100110001010101000011100100100101011000011001010101110010100011;
t_expected = 163'b1010010010111101111100001001001011000100101111100001000011000011101001110101011011111111010110001010100011111101101000000100011011110001111111001011101011000010001;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1110101000001100101011101011000011110001011101101011000110110001101101100111101001100000001011110100110011110101010011010101010011111101101001110011011111110010010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01100100101111100000000101000101111100010001100100100010110000111011011010000111011100100001111001000111000011100101101110111101001000111101101110011110101101100010;
t_expected = 163'b1011011001100110001110110010110010001101101001100101110110101001110110000110111100101000100010110000011110101010110001000110110001000100110001000110111101110110100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1101011010110100111110010111110101011000001100000010100011100011110110110011011111111010100010011001111001011111101101011001101100001100111011110101000001001000000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01011110111011111110011101110100110000001010100101111110110101111111111101000110100011010111011001011110001101011011100000110100100100101000110011000000111010100101;
t_expected = 163'b0000011011010000101101111101110101011101010101100001011100101111001000101011011110100110100001010100000001101100000111101111101010101011010010010010110001101110101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1111010000011101000111000011101101001110101001010011100000101101100001110101001101000001011111001101001100110110000100110000011111000100000001110010100101000010110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00100101000111110010000000011000110000111010010111011101001101100101100001001111010010101111111100010000100111001111100111101000100101001100001101000111000101110101;
t_expected = 163'b0101101001100011000000111011100001001010101011101011110000111110111111111000101110100011010101011100110100111101001000110100111000011110011000011110111111101010010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0100101011101110101010101100011001110010101010011110010001100100111010100011111011001011110100010011001000111100101010011110110000100000111011100000111011010000000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01101111010101111110101010011010111100100001100101110100011011110111000010101100001110001100110101101001001101101010001011010001011000101001010000011000010110111110;
t_expected = 163'b0101110111101010001000011011111010110001011100111100100010010010101011000000001110110001101111011010000001010000111110110100110010011010000011000100000001100101110;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0101001011010111110101010000110111010110011010110111110110100110000001110110001101110001000100101111100000000100000110010010101111011010000100101110000101101010010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00010100001000100100110110101010110100110010100100101100010111000111101101100000111011110100010000110001010011010110000100011001110100001000100111010010101001101110;
t_expected = 163'b1111001010011000000001100111110000100101100000111010001111101101101011001011100001000001111000000101100001101101111100000010000011010100001011100011110101010110001;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1111010001110011000000100100001111101001011111110110010101011100001100100000001001001010101101111011110101001111011000101111001000110111010100101010111011100001100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00101110010110101001010010100100110110100101010110001111000111011001110000101001000000001110110110111110110001000010100010000000111101101100111010010101110110101001;
t_expected = 163'b1001110100011000010111001111111101110101100010010101010010101010111011010111001001001011000000010101111101010100011011101010111000010100100111100111101011001101101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1100111011001010111000001001011011001001111110101111110001011100010111110110111111000000010100110110010001100111110001000111110101110111101110101100110111110011110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01110101000110110101001000010100111010011110111110110111101011011001010010011000110100101001010111000111011101110001101101001101010000001001000101001010000001101000;
t_expected = 163'b1111000110101100100101111011110110101100100101000100110111010011101110111010100000101010101110100011101111000101010100101001111001101101000100101000100110010111111;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1110001100011011100101010001100001111111101111101101001010010111001100101000001001111010110001001000011000101011011111000011011110011011010100011011001101001001000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00001111111010011111010101010000110010001101101101110110111111001011011111010001001101010001110010011101010111101101000001110101111100101101111000000100011110111010;
t_expected = 163'b0111110111101011100100111100110101010011010011000100011010101010100101010011010001111101100010111010000110011100100010111101010100001100001000011100011100001111100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0101000100100010010000100111011101010011001010000000101011011001010010111100011011100000001000011000101100000000100011101101001001101010111110011101010010001011110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00100100100000011011111011111010110110010110011101011111100111010101101000110000111010100011010011000100101100011001000110100100110101111010100110111111001001110011;
t_expected = 163'b1000100011010101101000011000100110001000000001101101010000001101011101011010100100101010001010001101010110011010010111111110111000000011000011101111001001010111110;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0100111110000010101101001011001001100110001001001001001100001011001001101010111101001011100001000100100000101000001101000000100110100100101101011011111110010001100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01111110110101000111100011101010111110100001111110001101100001000101000010111000001111011010100101101010100010100100101000101100010000010111010111111000100100110100;
t_expected = 163'b1111111010000011010000011010011001110111001111011011111111001111111111010011000100101000111010110011010011101010101101000101101010111001101010100110110001101010000;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1110011100111111100110110110110011001100111001011000001111100011110110111100000010010001011000110000000101100011100101001000011001001100010011001101000000101010000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00000111101011001100001111000111110011110010101110100000111001111111001111111101110111110000100100110011000000110010100101110101111101110111001000100110110011100100;
t_expected = 163'b0100000101011101110110110111110111101011000101110000001010000001000001010011011110111100011111001000000110001110111111101000001010000011100100111001011001101010101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1101000110001110011011100010000110111000110100010001101110100000101111101010010100101011111001111110010101001011100010100100101110111000101001001011010110101000110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01111101010011000000010101010101110011101011001100000001001101101101111000010100000000000100001001101010101010000110000011111000100001010010110111101001001000100111;
t_expected = 163'b1110100011101111100100010111001110001000001110110101000011001011000110111100011001001010001100011101001100101010000001000011101000101011100110100101100011110011000;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1110101111100111101110001100111010010110010101110000011000101010100100101010100010110001000100100011011001000001011100001000100111110001010001000111111010010010100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01100110000101011100101000110001111111001000111101011011000001101001110001011101111101111110101000100000100100111010001100000000001010110111101010101010011111110100;
t_expected = 163'b1000110001011100000010001111010011000101101011010000011001101001001110010010101010010100110001011111010101000111011000111101110111010101001100110111110101111001010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0110011101010111110011110001100000100011000100111100110001111110111011111101110110011010001111010111111100101000110000010101011000010111000011000000000100011000010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00001100011001010010100100111011110111010011101111111010010001110011011111011100011101011111001100011101011110101011100000001001100111010011011101110100000000110100;
t_expected = 163'b0011000011000100010011001000101000110010010111011010010011110100000010001001111000100010011101101111011001110010000010111001100001100000011000110101000011010100111;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0101010011101110001010000101010100000101100101111101010110110100100000101011010000000010111110001011100100110000011010110111110110101111111000010110011010001010100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01110111001000111010111110001011011101000100000101100010001111100001101000100100100010100101101011000111111000011111100110010001101011100110100001111011111111111011;
t_expected = 163'b1011101110001000111110110001001110011100000100011101111000001000111111101010100101011010011010010101101000100101000100001101000010100000110101001011101100111101110;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1111101001101011111111101001101000111101100011000100110101011111111111111111100010111000010111011101000001011010100111011011000001000111000110010000100100110001110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01001100010110100101010010100111011001011111010100001001001111010101100001100101010111011001001010011110110010100001101001001100001010000110111110100100101000101010;
t_expected = 163'b0011100010110001010010110100100000101001101010111010101001100001101110100111010001001100011000110011011000010101101010010100011110001011000100111110111010000101010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1100001010010011110000110100011010011000100010001111010100011101000100101001110100010010101110110001010101110011101001010110001110000010110100010010101000111011000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00010110101010100001001110110101010001101100110110101000110011001111000111101110101110101010001111110011011000110100000001001101000111000011000011100110010111101000;
t_expected = 163'b1000001001101011010001110010010000101101111001101100010101000111011101000110000000001100011101101100101010101000010101100101101100001010100111011111010101100001011;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1111010010100000001000000010000110100110010011001110100011000101011111111111000010001001010111101101111101111001000101111010110001101010101110000100010111101001010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01101101111000101001110101010001011101111111000111110000110111001111011010001011011000000010101111101001100110000000000110110101101011100100010100111001000000101001;
t_expected = 163'b1100101100111010111010111010110100111100001011110101001011101100011000111111110111011010101000011011011001111110110100111100010011110101100100110011010000010110010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0111111000011001110101101110111110000010010110000011100011000011010011101001100100110011110010111000111000010000101111010010010000011100010100000011101001010011100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00010111100100110111111001011001011101100100010101010011101111011001110001000011100101110000010000110000101100111100101000111110000010000000111001110110111111111110;
t_expected = 163'b1001100100000011010011001100001100001000111100000000000101100000101011000010010100110100010001101100100101100111100010011000100010110110100011001000110000001010010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0100001010111000100000010011001000111000110111110010001000001001001000111101111010111001001011000110000100011010010011011100101111010100111101000111100001011001010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00011100111000111010100001101010010001010000110101101010111011000011010110001010010100001001110001111010001110101111100101100011011111100101100110110000101100110110;
t_expected = 163'b1010001101110011110011010011000100010010101011100011110011101111101111000000011100100010101010000110011101000001101101001010110001110101101000011111011110100001010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1110000000000100011101000111010100001101100111111010101111101000010011101011001100000010100010010010000100110110111100110001110000110001001111001001010111001010000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01100110001011110010001111101110011000001011000110101110010101010011001010101011101010111111010101000111100000010011000011101011110011000000011000001011110011100101;
t_expected = 163'b0010001000101110010001010110110110101010010111110000000100101000110011000001000010111011010011010000111100000111000100000001001011100001011000100010011001001000101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1101111001111101100100101011100100101001000000111011011110110010001100111101111000011000010011011110100001011111010000001101010111001001010001011111001001110000100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00011101010111001100010011010100011000011000000010000101000101101001101001100010011011010111110100011100111010100111001100010010011010110000101101000100001100100100;
t_expected = 163'b1111011110101010111010100110111101000001100100000100101001000011001010001000111101100000010110010111111010011010100010011111000110001010101101111011011001001011000;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1110011111011100100011010101011010010111001001110110111101111000110111011000101010100010111010100010111101010101001010001101101000000111101011011001100101111010010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00000011001101000000101011010100010110001011111000010101011001111111100100100011100110101100010001000100010100110010100000001010011111010101110010010010011011100010;
t_expected = 163'b0101111001010111011000000001001111101010101111000011111000000111110100011000010000111110011001101111111111101000100001000001111000000100011011111010110010100111101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0110000101100101011110100000100110110011111000001111011001111010100000001110001100101000000101110100011110101101100110100001000011100110010001011110011011001000000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01111000011001001000100100111000011110110100001011111100011001111111011010011011010001011110010110101001011110001100100111000011110011111001001111011101100100110011;
t_expected = 163'b0000110011000001101100101000110010010100011110001010101011100010111100101110110111001001111111111110100101100010110000111111010000011110011001100110101101111010101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0001101111110101100011001100110110001000111101001110111010110111101001011000111010010011101100101001010010100110001000001100010110001010100011011000000101010010110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00010010000111010111011000101010010010100111001011000111000101100101011001010110101001110110110110110011111100111000001001011110011010111100010000000110110011110000;
t_expected = 163'b0110100111110000100111111010100111100010100101011100011010101100000001000000011100100101101111001000110010001101000110110110111011000001100101100011100110000100010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1011011110011000111010010000001000101100011101000111011101000101110010001110101100001001011101011101100110001110100101000010111001011010111010001100111001010000100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01001001110110010011001010001110010010111100111000000111110011110001110100010111011100000001010011101010000010101100000110011110010111011001100101001001001100111000;
t_expected = 163'b0101000000001010010111000000000110111010111001010111000110100110011101000110101101000100101111000111111100100111001000101010010011100111101101100111110111101001000;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1000010100101001001111100111111000010000001100100101100100001111101101011010011010100011010100010001100011000101011111101010000110110110000000001010110110101011010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01110011101010001111000110010110001110011111111000101110111011100011000011111110100011111001111010100000001000010101100010100111101011111101111011001111011001101111;
t_expected = 163'b1010000011010001110110101110101010011001001100101100001000110001011111011110010000101000011100001011010111101001011010101010001011110111011000111100011001110001100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1011101110010001110010001011000100110110101111101000100111000111110110001100011100111001101101001111011011101101010011000111100001011101111110101100001000100001100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00001000110100000101111110110100000110000100001010111101101111011001001011111111010011000011011101011101100010100001101101101111000010001110000110010000010010101110;
t_expected = 163'b0100100101000001010100100001001011111000001101001111011011100110100001010000001101011111101010000100001001010011101111110011001010000011111100010101001001010111001;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0011001100100000101000110111011010100111101010111001000010000100001001011010101000000010001000111011011111000101111101011011111110101101001100110110110110110011110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01010010100100101001110001010001000010010001111011010101100110011001100100110101111110100010101101000110001100111111100011110010000111101010111001011011100101111100;
t_expected = 163'b0000011101110001011001101000001111100010101000011111000101111011111010011011000100010100011110001000111110101100110100010010011001001101101010001101110111001100101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0000010010001001000101100110101010001001011011110000100000011010010011001100010010101000110001100110110010001110001000110111000100100001000110110001110010001001000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01111001111010110100001101001011001010100010111001100000110010000111110011010100001001011100101000001110011110001010000110101011101011001111101100001101111010111111;
t_expected = 163'b0010000111010110011011100011010111001111100011000011110000101000000011100001010001110100011010111100011000101000110010001010011010001010001010011111001101111101011;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1010111011111100110000001010010100111101011010011001000011111000001000011000000100110000011000100000100010100110100010010101100001000001111101110111001100000011110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00000011000111111110010101101111000011111001001001101000001110010101011011011001110000101100001001110111110000111110001000000011000010101010010011000010000101110010;
t_expected = 163'b1100001111000101111110010011100001100111100011101110010011000101100101101001011100010001011100000110111011100011000011001011101111001111011111110010001000010001001;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1001001001000110101101110100100000010001111110011000110110110000000101011111110010001010100001011000000111101100001110011000011110101110000111110001010110010100100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01011000010111110010111011110111000101101010100010001011001100000101110100000000000100000111101100101001011010100010100110011010001111001110001100011101010010100000;
t_expected = 163'b0010010010001011010001000100010100101001111000110011101010000001101111100100111001100101011100110110011111101011110000110100111001000111101101101001101010110001101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1010000011000111010100000001111000100010101101000101011101110011011110001001010100001001000000000100001011010101100000110100010001110110110011100101111010101110000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00100010001001101100100111010101001101110101110010110010010000111011100001100000111111110111001010110000010000000101100011010010100011001011110001110011101101100001;
t_expected = 163'b1111011110000101110111010100010011001001010111110100010111010111010110110101100110111111110111010101001100110110110011011000001110001010111110110100010010101001010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0010111001111110100001101101000111001110001100000101111000101001000101011101000010110011111011010000111011011011111110011000101110010010001001100011000100100100010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00011011010101101100101110010001000001000110000001110010000000101001001010101001001010001101101011111011100110110101001101000111101010111010100111110000111010100010;
t_expected = 163'b1100111100011101001101011000011100101011010110011100101001001001001111111011001010001010010000001100011011011011010111010111011101110000101000110101100110110111101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0001010000001111111110110001100111111000000001101100011011100001111010001011110100101001010110101110110110110010010111010000001101111010010011100100011010010110100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01100001100111100001010000101001100001011101100011001001101100101001001100101000110110110000000110000111001100101001000010011110010101011110011010101111100101110110;
t_expected = 163'b1001010111010001001000001111010011110011111000110101000010001011000001111001011100010010101100111101010111010000010100010000011111000001111001101111011010110101101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1011000010110011010011000101111011010100110000101101001001000111100001010101000010010011101111101011010010011010111001111101110010101111101000110010100111001100010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00101010111011011111001000101111101101001110110011000000111000110111110001000001000111010010000111011110000110011101100110110110110001111011100101100001010110110101;
t_expected = 163'b0010010010101110110010010111001000000011010001110110011100100111100000100011001100001100111001110011101111101110100110100010011101001111000110101111010101000010011;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1000101000010010001010101010001101100001110000110110101100001101111110000011010011011000001110110111000010010000000101000011111111000101011010111100001001000111000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00010000101100010111100100010111100101111111010000100000100000100111011010000000111000101010100001010100101000101000101001101111111000010101111000110110001001101101;
t_expected = 163'b0000100011101110010000000011011000001100010011010000011110000101110010101110011010000010001100000001111001111100001001011000010100101000010010001100010010110001011;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1001000110101011111111010110110101000011010101011011001111001110100101010111110101100010110111001011101111111001101011000111001000101001100000111010010111110101110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01101011110100011011111010010100101001100001000000011011100110110101011111001100001101011001010000101101110010110110000111100011010101110000000111111101110110101110;
t_expected = 163'b0111110111100100001110001110010000110000111110110110010001010110001010000110101001100110111000011001110111011001101100110010101010011001000110110100111110101010010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0011010110011010000010000010001001111111000110011010101110010110101100000001000011111000001110011101101011110011000010101110110111001001111110111100101001101101000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00110001101000000101110011110000101001110010110010011011111010001111100001100101110101100011110101110010010100000010010010111010111001010001010010100011100001101111;
t_expected = 163'b1110010010100010010000000101010111101000010100011100000111011000111101010110110111011110011001011010000100011001100010010111111010111111001010101100010001000000011;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0000111101110010011010101111011111001001000111010010000001010100110011010110011101010011101011000001010010011011001100000010011100010100001110101000101101100111010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01001010011010001000001111101000100001101001011011100110001010001011100010100100000010001111010101101010111110011011111100110011110000110101101000101100011110111001;
t_expected = 163'b0011000100100100010110001001000100100011011101101000110011011101000100010000111111101010010010111100000001010001110100111001010111110001011011001111110000010011111;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0010000111000111101101010001100111100100100010010011110010111010001001000010101011001101110010100101010110011000110000001110001011110110100100101011010011010101100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01100000000110000000010001001010101110011010001001100101000110010001001111011101110111111100110000000001110100101111110011001011011101100000110111101011001001111000;
t_expected = 163'b0101000100101011010101010010100100110111101111110110011110100001011010000111001000110010101011001011111010100010010101111011001110001110001100000000111010001011001;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1001000101011110010000100101010011010100110010101010010010110001010110000100101101110111011011111000000010100000011110100000100100011110011111101101101101001110010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00111011011001010110111001111110101110011001101001001101010110000011010001011110001111000100010111011001001010011001111111010110111000000101001010110001010110111011;
t_expected = 163'b0011001111100000010101111111000010001011010010111010110010100110110000111010011000010001000011011010110000010011001010101000100001000000111111110101100101101000111;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1000111111110110011101001000101001111010010011101111110101100001000101010010011011011101100010100110101011001011110110001001011001000011000101111011100001000100000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01000001001001111010100111110110100010000110011010111100011000010111110000010110111000100110011110000100100000000100011000010111100000100001111101111110100001100011;
t_expected = 163'b1101101100110111101100110001111010001000011010000111100000101110011101000010000011000010001101011110001110010100110100111111111101010111001100101100111000000100001;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0010010110000111100100010100110101001111010010100110110100101011011110000100101001000110000001010010101111000011001001010101111110100011110011111101011011110110110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01111010110101110011001110010000101010110101001010110111001100001100011111110111010001011011111010001111100010110000010110001111001101000100100000101001111010100100;
t_expected = 163'b0000000001001010000011110101100111001101001011000100010111101000100111101111100111010100001011011110000100100100111011001011110000100001110010011011010100000110100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0001000100111110010001100000000001101001100101101111010011001001010011010000111101111100111100001110011011101011000101111001100000001111001001110011000100111100110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00100000101011101101010010001000101110101100101001001111110100111100001000111010000100100001011011110111001100000100111001100110100000100100011111100111000111110111;
t_expected = 163'b0100100001011001011111101111011010001100001010010111001000010001001001001110001010011011110010100000010000111000000110101110000101110001011100011111000110000001000;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0011101010001001001100001111111011010101101100011110101000000100001000000110001011100110010101001010010110100000101011011100001011001101110001110110111000001110000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01001011111011100001000100101010100110111111011011101110110000111110100000110011111010010001111100101000110110011010111101111110101000000011000011011100000000110111;
t_expected = 163'b1000000100100110001010110110100101011001011110100000110110001100011110011001011001111100010011111001010010011101101100101011101010001110110110111011101101011001000;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1000010000100001110011110011100111110101001100010000001000011110110011010000101101001110100100110101110100001100000011010100111100110000101010100000010110010100110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00110001100100111001101100111111101110000000011011100100100000100000101111010011001011111010011101110000111000101011010011110001000101110110110100010011111111110100;
t_expected = 163'b1001000110100000010010110001010111111000000101110001100010101110100011000010011000100011000111111110101010010110100010011110111110000101001000110100101110100101010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1001010000010000000010100111010011001010011001010001101111011100101100000100111011010101001101101001101001000110110100111010000011011000011000000110001000011111100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00101010110000110111110000010111100010010011100000010101111100110000011010011010110110001010101001011011010010010111011100101000101000110010101001010101101000101001;
t_expected = 163'b1001011100001111000000001101101001101010110101101101011001001111111101110001101101101000110011000111011111101001011010001001001101011000011101001000010011101010010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0011101011101001001111001011101001101110111000111000001110010110110111010011000101101111110100111101001101101111011000010110001110011100100010000000111100101101010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01010000001010111010011011010001100010000000110000011000011010101010110000001011000000110100101000000010110000000011111000110000101000010111010110001010110111101011;
t_expected = 163'b0111000111000001101100000011110001001111101101011101110111001011101010000000101000101111000111010110000011101110011100010110110100011011101111010010010001010111010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0000000001101000110010110110011101010000111001101001111101110111101000000101110011100101011101000001001101000101110110011011111001100110011100000110110010110111100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00101011010110000100000111100001101100011011010010101010000010011100111111100010111001000101001101011110101110110110110111011001010101110010101001000001000000101010;
t_expected = 163'b1010010000100101101101010101100110000111010100000010101001010001100110111010011000000100111001010100011101011001001101000110100101000000100111000010100111101000010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0010010011010100001110000100000101110000001110100000011010101101110010010011110001011111101000000111110000011100101110110011010010000011000110010000001100111101110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00000001000010000100111011101001100101101000100011000011010110001100001010101111001100101111100010010101000101001000011001001101011000011010111100010111011111111001;
t_expected = 163'b0001111110101100011011001011101110111101011110111011001000011101110110001011010111010011001011101000011101101011011111110101011111010010011101010001101000011110101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1001111011100101011111101000111011000101001110101101011011101011111011010111000101000100000001011011110100110100000000001111101101101011100101010111110010001111000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01011010011000001000110001011111100001110111110001000011011010000110000001101111110011010111000010101101001111011100011100000100110100111111000010011000101100111101;
t_expected = 163'b0100000111010010100010010101110001101110110101111110011101110001101100000110101000101011000100110111010100111101110011010011101000000111100011111001101011110110101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1000000101001100100000110101001111101011101111001101110101100011000100000001110011101110111000100110011100111110101111000001100010100111011101011111111110010100010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00100001000101010110101101010111101001100100010000111010001010010000100101000110000011100100100111110110101001101101110010011101011101011011011111000111110011101110;
t_expected = 163'b0010000111001001010010110110111111101001111111100001011010111011111010101000001011110000110101000000110011010100111101100100110011101101010100011010010111111111100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0010000110111100011101000001110111111111111010000100010100101001011111010111100101110100111011110010001001010111000011100100010101010111100111001001000001011110100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01011011100111011111000000110001000101010101100010110001100100000000011010000101111110001000000110111010010011010001111101100101010000101110110000000101001100100111;
t_expected = 163'b0010001111001111110100000100100100111001100110111010010011011011001000101100011000010010010010110110010001001111100110110010100110001011111010001111110110100011010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0001111100000101011100101111100000010001011011010101100111011010000000000001010011001110000010101100101101011101111001001100111000111100111001001111111111101100010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01000000111011010011011010000001000101001111100010000001110100011010010001001100001001111010100001000011011001000111111001101100110100001011100101001010011011100101;
t_expected = 163'b1101010010011000101100100111110110000001011101000000000100010000000101100011110010010110011101110110110110011110000100001011010101011010111101010110010010111001001;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0011010110110000100001010010011100100000011010011110000000010000011011010101010101100101101111001100110100110101110101000000000011111000001011001001100111110110010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00111010101111001101100110001000001101011100011001101000101000101010110101101101110001000001100001011000110111110010010110110000011101001001011010010101000100110000;
t_expected = 163'b1001110111110010001010110100111001101110010100001100111001000001101110111101101010001001110101111000110011000101110111101001000100000011011110010100100010000100111;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1000000110011001011100100110100100011100100001111011100001010100000000000011100111111111010110010000010000011110011011101101010100000000110000001110001001011100100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01010011110101000101101110111110000001010011101011101011101101101100101010110101000100111001010100000100011101001110011100111001010000101100100111011011110011110011;
t_expected = 163'b0000010111110100010101011111111010001000000001010100010101010001110011001000001000011001111100001101101100110100010011010000000101111110000001011100001000101010011;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1001101101101001000001101010110010111010100101110010000010011110001101010100010001000101110111001100011100010110100110000001111011101101001010011000011111001111010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01001001001000101001110000111110000001100000101011010111110101110110001011111000111111011111110101001111001011011010111001100000101110001001111001101000101100110011;
t_expected = 163'b1010001101100101100001111010010010100001011110100100100011001011101110011011000000001100001000001111101111100000000111110010001111101100101001110110000111010111100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0011010111110000110010010110001110001110000100101010111110001101110110000000001111011110001110111011101101111111001100011011000100101101011000011110100011000101000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00110010011110111110001100010110001111111011011000110110000001100110000100011001011010100110011001110111100001100110110111001000000111101101001100100111011011101000;
t_expected = 163'b0110000101100110111110100110111110110011110110111000011111001000011100101110101110000110001001011101111111110011111111110001110110100011100010111001000000101000011;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0000010101010001001111100001111110100101010101001011111101100101101101010110111011110100100111110111101001100001100000110111100011010011100000011010001101111111110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01001000000110110110000111000000000111101000011000101100001011111000111010010000100110010100111110101100001011000101011000011101001010011000010011111001000000101101;
t_expected = 163'b0111110110111101110111110001101000011001010100110110100010100101011110110111101101100111111100100011010011000010101011101100000001001011111011110101100111001101010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0010101001101110010010001101000000010001110000000010011010101111110010000000011101101110010110100011000101001001001110011010111111110011011110000100010011101101100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01010011011000111010111011101000001010011111101011001101011111001010011011010001010101111100011111100001000101010001011100000101100110111100101100111110111111111111;
t_expected = 163'b1000011100100110111111100100010010110101100101000111110110001001100110110110101101010010110110000001101011001010110100101000000101011101011101111000111111101111111;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1011000011010110110110010001011000111101110001000111111011101001101000000110001011010100101011011101010000000010010011011110010100011110110100000010101100100111010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00111001001100100100110111111110001010000110011011000100000011011010010100111001101000000111011010011001111101101101110010001100000111011101110001110101101010111100;
t_expected = 163'b1110011101010111010001100100100111000000101011111000001010100100001000010110100010010100011100110101101110111011110101000001101100101001100001011101101011100001110;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1000010000110111001111100100101100001011100011011110011000110010110111010010111100011111000010000001111000101010111001110110100011010110100111000101100000010101100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01000010110101101000001101011110000010010101011001110110100011010000100000111000011100110011111010000010011111011000111101010101001010111000001110101010110101111101;
t_expected = 163'b1010011000100000000101110011011011011011000001111100101001001010100110001100111001000010000100100010111100010000010100000110110111100000100000101001111101010101110;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0010111010001110010010001000000010100010000110110111101100110010100100000100001110100111111001010100111101000000010101011000001100100000011101000011011110001110110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00011000101011100001010001010110001110001110100000011111111111000100101011110001100111001001011101011110010001001110011011111001100110110100111010100100010010101111;
t_expected = 163'b0101101110000111001110100010110010101000101010111010010010000111000100101011010001000011100010000101100010000101101111110111101011011011010010110110011111110000001;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0101000010111111101101110110110010010100000111110110000111011000001101011010001000111101011000111000001001001001111011010101010011001000100111010001100000000100000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00100011111111011111011000100001001110111101000010000110111101010110000100011100010010101001111100010101111011110010010110100000101111010011100101110011001101100010;
t_expected = 163'b1001001101011101110010101101011110010101100001111101010111010110000001001010100110111011111000110100001100111101000010010001101000100010000011000100001110011111100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0111000000000011011100000011101110110000110110111100100100010010010010001110111110010111100001101110000001100001000111111001100100001101011111010101101100110110110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01011001100101010011100110101001000010100010010010100100100001001100110001001100101111010010010001101100100101000011111000101001010010100110011000111000111010100001;
t_expected = 163'b1111111011100101111101110101111100110000010001100010111111110010111001000010010001100011100111001111001101011101010111101101001011000100110110001100001000010011010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1110111011000010000001011111010000001100110011111001000001000011001001011001001000001100001100110010110100101010000100000001001101110101001001010011011010101100110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00010010010001000001100010011101001010110001100001101101110101111000111011000111011111100010100001110110000111011111111111110001111110000010000111100110100101110001;
t_expected = 163'b1110100000000011100001000000101011001011100100111101010110000100101000111000111110111101110101100001010111010101000001101110100100001100101001011110110011111010101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1101010101111011101100110011100000101011010011000000100010001101010010001111011100110110010101001110111000000010101000001100110010011101110010100100000000000110000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00101000001101001100011010111111001100000010000011011001011101111010010110100110100000011100000110111011101101101011110011000000111111100011110010100001010110110010;
t_expected = 163'b1001010111010010010011111001100000010101010011100110000110100010110010101001000001101101101110110100011011110110011010100101010010101110111111111111101001111101111;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0111000111001011011001000100111100010011001000000001110011001111001101011001100010001100110100011010111000101000010110101000110101011011001000101010111100010101110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01010011010110000000000100110111000100011001010010110010001001100000000001101111010001110101000011000011100011011101011100001100010010000111101101101110001001100110;
t_expected = 163'b0110011111101101000000101111100101100010101110011101110010111010001100001010010011101010101011000011100100100111011110111010100101111111101000100011001001100101100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0100101111100010000000111000001110110101101101001000010101100101010110001101100100000110001101010101001111110001111010000110001010110010110010101100010010001111100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00101001000010011010101001000001001000001000110000110011010101110100101011000110101101000111100010011000011001000000011010010101111110100010010111010100010110100101;
t_expected = 163'b0001011100101000011001101001111111001101110110100110010010100010001100001011010100001101101100101111011001010011100111111100000101111101001110101101111000011101001;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0110010101010111111111110100110010001000101100100001110110110101011011001011010110111101100100100001000011011011010001001110100101000110100000101010001101100101010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01110010011000010110110001000001000001110111000000001011010111101110001110000010011010111111000110000001110011110100110111011100110111000111101010011011100001101100;
t_expected = 163'b0111001011011010100110100001111010010111110101000011011001011000000010010011001000010110110001001101011011011100111001011010000101011011110010111010100100111011010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1111010110101110000010000000001110101100011101110101011011111110100000011101100000100111010001111101100010010111111101100011011010101110011110111100110011110111000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01001000100100111010111111111001000001110100011011101000001011111100010001001011100011011000100111101111110101100000111001000100011010000011111101001100111110111110;
t_expected = 163'b1011100100011111101010101010100001110101100000010101110100100000010010100111111010001111110011011100100100111110010000111001111101100101101010111110011000110110100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1100101100001110010110111001011100011110011101111100101000110000111010001001110110001101111000100001111110111110100011001111011011100001110111111000111111101101110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00100111110000100001000111111111001101100110111011110001111011001100111000101010000110100010000000110110011111011011011110111001110111110010000000000010001001111011;
t_expected = 163'b1010011100100010001010001010111001011011101010101100110101110101011101000101110110101000001111110101111111001000010110101001001011100111010010100000001011001110101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0110000100110111101111010111100000100010111000111101001001110000100101011111010000010111000011010111011010110100001101000011100100010001001101111111000001000110000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01111101101011101101011011010110100101111101101001011001110111000010111110110011110000011010101001101110100001101111010010110001101111010100011111011101010110111000;
t_expected = 163'b1111011011101001111011011101000111000001110011000001010001101000011100110001101001011111000000010111100111110010111110000010111110101110000011110001110100000011000;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0101010110100100000010100011010100000101101011010100101110001010111110001001100100100100101010011011011011011101100001111011011011111101011111111001111111010100010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01000110110111101001110100000010100001001010001000011010100011010010000001110010001001101001101101100001101011111011111101101010001010110001100010011110100001101000;
t_expected = 163'b0100001000010001011110101111011001000010111111001001111111000100110101010011110010011001101010111111001110001001111011110101111001111011100011000011011101000010101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0111111001011001010111111110101110111001001010000011001100001001100001011110110010101110011011001110100111110111011010010100111101111101100101101111111011011110100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00111100000001110111101100100000101001010001111010100010111011000000100100011010111100000001011100011000000001000110111011100011100111010100110100000000111010100011;
t_expected = 163'b0010100000111000101110000101000111001011010110110001101001010000011100011011101001010100001010000000101110011011011110100000000110010100111100101100111100111101011;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1110000011111001101100010010110011011101001111001010001101000011111010001010000100010100110010110010100011111111110110010000100010010000011111100101000101100100010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01100111011001111111100010111000100111000010101010000111011101011110101111010011000010110111111011000010100111110000010111110011101111110000001001001111100101110100;
t_expected = 163'b1011000001010101001110011111101010110011100111000011111100101000110100001101100111010111001011000101111000010110011011000001001101011000111011000001111000011001100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1101001011000000010001100100000011100111101111000011110010000111010011011100110110001111001111101100000010010100111000111100001001101010100001100011111011110110010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00001101001111110010011110011110100111111001001001011110000101101110010011010110110011001110011110001011111101101100011000011110000010011101110110000000010010110100;
t_expected = 163'b1101111101001111101011010101001100100010100010100010011001000111001010101000101010100000100000110011101110101111011011101000001111010010001001010110010110111010010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0111111001110001001100011001111101000010111110100011010011011101001100001010111000100101101110111100011110001100010100010101111100101110010010110100100111011101100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00110110010010001100000110011110101111101000111011111100000001100100010100111101001110100100111110110101010111011001111110000110101111101100101011010010001111110111;
t_expected = 163'b1110101001100001111001101100101101101101111100101101011111000100101001110100111000011011001001111001010000011111010011001011011011110000000001000110101001111000001;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0100010011011001111001010101101001010100010011101010110100110110010111011100001110111101010111010000111011100110101111011001010011000110001010110000001100000111110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01101110001010000100101001100010100011111111111010110101011101110110111111111101111000010100011011101100011001101001110011011111100101101000011100011101111000100110;
t_expected = 163'b0110001000100100100100000011110110011111000101001110010110101111100100001011010000000100000111000111100110101101001000001001111101001110010110101110001101101010010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0100001000101100010000100001010001111000010000111111010111110110001100011000111000000111011110000100100111101111000011110111001100110111110000110110010010010101000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00010101111100001000110001100000101010100100000000000100001101100010101011110100000001001111111010110100110011110101011101010110010000001101000011000010100111100000;
t_expected = 163'b1111000101111011101011000000101011000101011100010100001000111100010001101011101111000001001111000110100100000111111101110001000100101100001100011010001001111001011;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1111101010010101001101011100101111001000100001010110110111111100010011001110101110111100100111011011000111000111101101001011101011111001000010110000101110111111110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00101111100000010110011101011000101110010111110000101110100011111000000100010101110100011011110100110111000101000011011010101010011101101001111111000100000000101001;
t_expected = 163'b0000101011010100000011100111010000010101101111000100000000010100001011010011010111000010111010110010000011100001101000001010001100010101101001011011011010101100001;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1100010010111100111010110010011011100111100100010111000000111110000000011000001010110110010010100111000010101100010001000010010000010001111100100110000000101101100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01100100111010011111000011111101100110001100110011111111110111101000101101001100001111010001010101001010001111110110010100100011110101001100100000111111011111111010;
t_expected = 163'b0111010101001111000110111100100110010110101111000110000010011001011111001111000010100000010100100111100000100010100101000000011011010100011111100000011010011000110;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0110011100101100000110000110000011010011000100011110100001100000101100001100011100001100111001100011111110100100011011101110101111110101110111100000011110110111010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00011110101110011001011011111111101010011011000011010111101110011110111010000101111011100000110000010000100101101010111001111011011000101011010101110000000100111010;
t_expected = 163'b1010111100000000110110110110000101011011110010010010000000000101000011100110000001101010101000011000111011110010000110110011100110011101110111111111111111001111101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0101111111010101011111011010111101111101010101000100101010001001110111011011101110010110000000111111111110001010111110001010101010001100001101101111100000011100100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01100101110111000101110110000011101000101000000001111100101010010100010100100001000110011010010001011001001011011110110111111010010101001011101010110110110011101101;
t_expected = 163'b1111111101001110001101000000111101111101001101110100101111101001111100010111001001011101001101101100001101110110110101000011100001111110000011000000000111101011011;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0101000101100100100010110111001101001001010100100001001101001011101100001101011000111101100001000001010011001011010000000110010101001000111101111011100100001110110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01011111001001101001101000000001100100100011110000101101010010000100010101101000010101100110100111100111011001101101010000100111111101111110110111101001101100101100;
t_expected = 163'b0110110010000011011101011111110011110011001100110010010111001000110010111101010010001100100010011000010000001010100101011001011011001111101001110111001101100111000;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1110001101001001000111000011110001100000110011101000111101000001110011011011001110100111011000010100000111100001101100101101111010100010000111011101011010010100000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00000100011101110011001000111001101100110010000010000001000110010010101010101001101001000101000010111110110011110001011100011111010000111011001000100010011011100110;
t_expected = 163'b0001101110101010010110011000101000011011011011111010101101000000001000001011110110110110000101101101001110100101101110011110100000001011110100100111111001101110000;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1101111111111001011010111101100111010110100010101001011110010001101000001111100000011001110101001000100110111001000110000001101101011111011101011011100100111110010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01101110000111111110010100111101101100001001000011010010001000001000000110000000001100111111000011100111011101010101110011010110010101011111010100111100000100110111;
t_expected = 163'b0011100111001010001111011100000011011001000111011101111100000000100011100110000111000110011001111101001001010000010101011011100001000011000000110011011000111101100;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b1111010101000010100001110000011111110010000010100000111011011110110111011001010111010011001100101100101010010000101010001101000110011111100010011001111001101100110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01010101010011110010001110011111100000011110111001111011011000011000000101000001110111001111100110101101010111101000110101001111101001111010100011111011110011110100;
t_expected = 163'b0111100100110000101111010000101111001001100100011010010000101000100100101010111010101001110011110011000111001000000111010101001111100001011000101001001001110101010;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0100001110100011010100000100100011001100000111010001011000111100001100001111000011101000101101110010011110111010110101110000111001110011010000001110010111010111000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b00001111101100101000100011000111101000000100011011011011010100110010111010001001000010100100001110010000101001111100011000000111000000011110101100100100101100110000;
t_expected = 163'b1010110001011001100100110000101000110111100101100101001010101010010000010101110000010111110000010000100011110001101100100011101110110000111011010100100100000011101;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;
start = 1'b1;
a = 163'b0100101010011010001001111000110101101101111110011100110111110110000101001011110101110010010100101110010111110011011001011000010101010001101010001000001001011101010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 164'b01110100110100100100111101100010101101010111001010000000100100100100110111110110111110011000101001001010001011001010010110111010001101110111010001101110111011100011;
t_expected = 163'b0110011000010001101000101100100010101000010001001110101011001001101111011011110010011101010101001000101111010000110011110011100010000011011000110011111101011011000;
#20;
start = 1'b0;
b = b_total[163 : 160];
#20;
b = b_total[159 : 156];
#20;
b = b_total[155 : 152];
#20;
b = b_total[151 : 148];
#20;
b = b_total[147 : 144];
#20;
b = b_total[143 : 140];
#20;
b = b_total[139 : 136];
#20;
b = b_total[135 : 132];
#20;
b = b_total[131 : 128];
#20;
b = b_total[127 : 124];
#20;
b = b_total[123 : 120];
#20;
b = b_total[119 : 116];
#20;
b = b_total[115 : 112];
#20;
b = b_total[111 : 108];
#20;
b = b_total[107 : 104];
#20;
b = b_total[103 : 100];
#20;
b = b_total[99 : 96];
#20;
b = b_total[95 : 92];
#20;
b = b_total[91 : 88];
#20;
b = b_total[87 : 84];
#20;
b = b_total[83 : 80];
#20;
b = b_total[79 : 76];
#20;
b = b_total[75 : 72];
#20;
b = b_total[71 : 68];
#20;
b = b_total[67 : 64];
#20;
b = b_total[63 : 60];
#20;
b = b_total[59 : 56];
#20;
b = b_total[55 : 52];
#20;
b = b_total[51 : 48];
#20;
b = b_total[47 : 44];
#20;
b = b_total[43 : 40];
#20;
b = b_total[39 : 36];
#20;
b = b_total[35 : 32];
#20;
b = b_total[31 : 28];
#20;
b = b_total[27 : 24];
#20;
b = b_total[23 : 20];
#20;
b = b_total[19 : 16];
#20;
b = b_total[15 : 12];
#20;
b = b_total[11 : 8];
#20;
b = b_total[7 : 4];
#20;
b = b_total[3 : 0];
#20;

if (t_expected == t_i_j)
	$display("this data is right");
else
    $display("error, the data is not expected");
#20;

$finish;
end

endmodule

